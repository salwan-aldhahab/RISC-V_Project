/*
 * Module: alu
 *
 * Description: ALU implementation for execute stage.
 *
 * -------- REPLACE THIS FILE WITH THE MEMORY MODULE DEVELOPED IN PD3 -----------
 */
