module execute_tb;
endmodule : execute_tb