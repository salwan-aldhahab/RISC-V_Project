/*
 * Module: igen
 *
 * Description: Immediate value generator
 * -------- REPLACE THIS FILE WITH THE IGEN MODULE DEVELOPED IN PD2 -----------
 */
