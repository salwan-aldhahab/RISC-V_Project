`define MEM_DEPTH 1023
`define MEM_PATH "memory.hex"
`define LINE_COUNT 256