/*
 * Module: execute
 *
 * Description: ALU implementation for execute stage.
 *
 * -------- REPLACE THIS FILE WITH THE EXECUTE MODULE DEVELOPED IN PD3 -----------
 */
