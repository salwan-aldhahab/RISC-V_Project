module register_file_tb;
endmodule : register_file_tb