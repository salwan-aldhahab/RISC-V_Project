`include "constants.svh"

module control_tb;
endmodule : control_tb