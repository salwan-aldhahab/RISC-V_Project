// ----  Probes  ----
//`define PROBE_F_PC          // ?? 
//`define PROBE_F_INSN        // ?? 

//`define PROBE_D_PC          // ??
//`define PROBE_D_OPCODE      // ??
//`define PROBE_D_RD          // ??
//`define PROBE_D_FUNCT3      // ??
//`define PROBE_D_RS1         // ??
//`define PROBE_D_RS2         // ??
//`define PROBE_D_FUNCT7      // ??
//`define PROBE_D_IMM         // ??
//`define PROBE_D_SHAMT       // ??

//`define PROBE_R_WRITE_ENABLE      // ??
//`define PROBE_R_WRITE_DESTINATION // ??
//`define PROBE_R_WRITE_DATA        // ??
//`define PROBE_R_READ_RS1          // ??
//`define PROBE_R_READ_RS2          // ??
//`define PROBE_R_READ_RS1_DATA     // ??
//`define PROBE_R_READ_RS2_DATA     // ??

//`define PROBE_E_PC                // ??
//`define PROBE_E_ALU_RES           // ??
//`define PROBE_E_BR_TAKEN          // ??

//`define PROBE_M_PC                // ??
//`define PROBE_M_ADDRESS           // ??
//`define PROBE_M_SIZE_ENCODED      // ??
//`define PROBE_M_DATA              // ??

//`define PROBE_W_PC                // ??
//`define PROBE_W_ENABLE            // ??
//`define PROBE_W_DESTINATION       // ??
//`define PROBE_W_DATA              // ??

// ----  Probes  ----

// ----  Top module  ----
`define TOP_MODULE  pd4 
// ----  Top module  ----
