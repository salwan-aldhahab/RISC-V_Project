module branch_control_tb;
endmodule : branch_control_tb