module memory_tb;
endmodule : memory_tb