`include "constants.svh"

module decode_tb;
endmodule : decode_tb