// ----  Probes  ----
`define PROBE_ASSIGN_XOR_OP1 assign_xor_op1
`define PROBE_ASSIGN_XOR_OP2 assign_xor_op2
`define PROBE_ASSIGN_XOR_RES assign_xor_res

// Define other probes as required....
// `define PROBE_ALU_OP1 // ??
// `define PROBE_ALU_OP2 // ??
// `define PROBE_ALU_RES // ??
// `define PROBE_ALU_SEL // ??

// `define PROBE_REG_IN  // ??
// `define PROBE_REG_OUT // ??

// `define PROBE_TSP_OP1 // ??
// `define PROBE_TSP_OP2 // ??
// `define PROBE_TSP_RES // ??
// ----  Probes  ----

// ----  Top module  ----
`define TOP_MODULE  pd0
// ----  Top module  ----
